library verilog;
use verilog.vl_types.all;
entity SPKER_tb is
end SPKER_tb;
