library verilog;
use verilog.vl_types.all;
entity CNT138T_tb is
end CNT138T_tb;
